BZh91AY&SY��� +�߀py��o��?���`�}Y|=
 ]��pܐ w ���8��m 	 � ��((!
����4�d�LOQ�4@�4	*P�F�`#�dɓ��&	�F�!�j~E(�&�4 �F��@� 4��=L�z����Bi�0��C�L�41I FS)�m&�<������?Q=ՄPC�.�EBʂ��(��÷�ʠ�
�/I��x@T&D!DO�i���I%��GD�A�(O$�����l����~K�0����nU���ʱn����U�y�z�Ԗ#�*b_
�9�:�99�4�z�	͝��ՑȀH�3h�8�����`'Cw����&�a/����"�}�ͮ�]Mv]K(��{��y$�ӓ��i���Η��F�)�r�g@��IWBSm�<M�t�ݸ�2��gNn�-�H�U
�I�,"E��n�$Ҋ�.�D\�|D����INSn�c�����B����M�;N�k���+|p��a
�Β���v�KGn�D�ɻ���|u�a;ٍ� Ym�HA�N`�Cb�>�c���b��N6�ֶ�jlط��,�;8N���t�:�\�J�i�ޏ���bhw%�գ����n�wt���/Z=��ٞ��G�í�M�����we��޺�6�V
�䳸ٚ��i��M����G�Mc�:A��9��[(4�����Z�M�����=�c�w;�:�s4D� ·{׭��u-W��cUN���\Y"7K��t��d:uc7T-�|�^�w����wk�N�vL�m����a���'�*BD\�8%��9��eY��.f���
%�z�yh����"r�N&8�iE2���f"y=���v��7�/�4�xx��t�͔۔�X2�s\��;�Ap�B��nfY��w�R��6���f�4ڦ؍e�&���֭�R\��m���i��8x3f�[�	��H�������Rl0�Y��!p����m*�V��5���jr�%��X�XF ���l���P&A��{�u�3/mD@9
�\�o�C���n5?X�����K�܅�Q"��	H�"�DC*��ׂ !!	�׽opn���;��xA��V,6�%����6,!�Bq1�,)e� J!UCTL���L@�Y�r�!al�*D�@R0����Rro*M=�_G�|��|���ۙ��s���Ɩ�
��'4���&�9��M��#�<��-��AD�0�� �� ��}~"�� ��"z|�
Y>~�4D�@ �6px��[�{� �xI�I3�JfH[Oe��&uU@�N` �/@ }|��X��m�X�(������hc��u�!@x��r�7U!
�e������*&���6�{� .m����YA�5�&
�����tM`2" ���ɘ^)��3v��1Tl0fֈ�b�� ����>�C��&���0�"�!�o�wL�~�f����hȔ�J xT�Z��
1�|��>6�e�� ��ϥ���sF����V0DG5
h� #
���D.#|�h�@�pu��@`RP�L�CĔd)�x�`Dq�^U$������������[z�;tj�f ��X���:Ü�  c�" {��ő �1V�vL���qP�30,��"s�%�$Qs�$!���8�sl�xF�n�]H��%L.�q�����qe�X:�)�g��>�&f�g�]6��E"��܀�YCB{�GwX���������u���~�|ND}7���2f�ҨSϐ���� ;B*}#�3�o&�" x��U�FP�S�T���tJ�p4�vfi2�X)�2@ �t/���=V�EQ��=��� :�D����f"I�>1 G��n�n� b� YSq�wp��2����e��\zIA1��<��0H�>����q��(�H*�~�z�H��zZ��zA-�D@�J)[Z�˭ii{�x���y������ZjEv���'���Ɍw��X&a˖�v��M\������,�YyKr�F�
�|t�+s�f�\���/3SB���q(��R��$����$��t���^*oPID��.K6����3� @���z}��w���>3�?s�7�x?R�� F��ެ�-?  U����.+�y}�_.���A��ﭫ���!!�"@"�Ƣ@2Й�>�0n�ƀ3�A\��X�lM��[fi��M���Ԗ)�K�mرW�`w��Z��(�߇�����Fed�.�/���M�M��~x"ZG�B��PM7>�͜�Ç�+����6�md�c:Ȉ�E��0		�9g��1&L�KfhXe�f�Dq�1����Ѯ4��r���5�nk��A�C` =�r<lt?S�)$��,ů<��t�o '��Q���щr��d"&Z�(V��^Mx�ϕ)(�w��>X�T?,D@/�0�X�	�`���	DA0�$"=�=qv��S8� A� K=�DU�L1)�B��Wԫ��� u��n�^�3ՠw� ��|�H� ��_������j?!<�?kg27E�]k��*UU�� ��ڑֳ�>��=�����N�{#��Vo��,Ȗ�R�.�/<��o��X�Z)11I�d-��!�K�Z^@��i[�MWz�M?�z�����Q E��y��������U����� ��!��#�" ĉN0���RDa�Q��=	���k���h֓i�R6dP�YIc�9�Rl��H%�2 � ���c�RfU�5-yuPz�˥��>����xwV��BH������&ɷ��Бk~� 	�$�f99�5њ�F縀�����0I$���*Z2뼿h�3�wz� g/�k���1�&K��b��}1}\��~u���ƍ�N&��׬:�@����� @�#�~�ȑ~5&e�ʓM�WH�_6r0��k�GҬn�e�s~\hz����  E��V��o|X���8:5�U7R}CcI�����XI�A�4�!���uyi��R����Q��>��~5�f{ 8I01��� I �#!].b��{2�
�3c$�49�=�/|B�^e�}�|is����F�~���{�N��k��ެ5��K9��׻rcCN͚�=��0�?H^�?|MQ�.z�Ɯ#wn�ɓ8����K&�BH$D�p=sӏ�����#8Á#��`
 �D\k�$����7H,���L�pp�h�#��4�`�r��F]���BM��NN��oU~(Wŋ})l��s��?���^����#RU�g�mIK>?&<n �a���4`�E�8<ċ��՞�9��ُ�5�j"!�Dx�d�.i!���E���ìO
�W�ueu���CL�U|L��� �\;u�\8���J�/0@��U���T�3N�r�[��8��&��A-I� �T˿�����3<u�O|r�]Ѫ���#�����!(H�*1aW�DXF<���	p@U`����s�Ar3/�-��Sz}F�xH����wW���D�wه�É���x���@ �`~��UB5UG�i���a
@��8R8�" �^��O�e�ځ�.��<��ٛ�  Fg��@��c�C���}b1 
悒��i&�2�����ػ/�?�}O]�|��Nh���2滦�j���E������DDR�N���6ڴ%�uo;��	�>��$񄄒I$�,D(�� �w螔�!v��
m��lkd�����R�44��F����L�` �q*Ė%	yJ�	�K�@�Q(RJ�DJ��D**�Q�Da��7���J��oK#%DYA"�
�@Z���HD[�6�/�H��6�!�Ԍ$H�d$
��qF H��H$$ ��f�E�I c1MH��zHH��I$FID!{K�!# 2 ��*�$�@�R����U"B�*H�X��7C׭� 0 �=h��BAIBADtCj�68����>�]9���	�`�U�!��񍟤�W�:�6�M ��,zBR�@��uS�CQ��'��iRuP�S5��3�����H;�""�%J�A�67=�w��@<�`��t�PH�s�!��5{"m)��'4�	�H*QD�l����ʝga҈S�&�I�[�����E��_<D�g��ul)�H0	����|>�����4<Ap$�t5x� !���F3�F��?��y�>$�C���R���j�lH @�DH�� ��ă �F%*����� �
��#p L�%h�7���s!�޸J	��'��L�� �A����v08��*l���I8��@��}�9s�>G�W�?g�酫�у��Pf�e���'܇�'gr\����-	�ɔ_7i��0�y��L;�&��
���������4�
��@H	^���yn-�暚���w��B�8����dK������)2��1������fR�9��'*.<�I��2]��|@:�����1���V�h"ک i��?�)��h��ǒB���~���a�'d�M�;��q��P���ntN����Q� ]�㨵��M3&$&D�b%(�l��8�x�%�{a�I��Ј��Q�
�J���0�&��2PP�g'	 ĺ��C����F���!ޅ�=�7���K�۶�<�S8-�D�wc� !��'7�I*H=��b����M��Q(���ƔX0��J-H��HJ�) ��{3�K���DNh���c	�7��.��nY�z��c
)�}q�Q�-^�@�E�`���"�(Hsq 